`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:07:08 10/19/2015 
// Design Name: 
// Module Name:    Imem 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Imem(rdadd,out,reset);
input reset;
input [31:0] rdadd;
output [31:0] out;
reg [31:0] add;
reg [31:0] out;
reg [31:0] mem [0:64];
reg [10:0] k;
initial begin
	for(k=0;k<64;k=k+1)begin
		mem[k]=32'b0;
	end
	mem[0] = 32'b00100000000010000000000000100000; //addi  t0 0 32
	mem[1] = 32'b00100000000010010000000000110111; //addi  t1 0 55
	mem[2] = 32'b10101100000010010000000000000000; //sw t1  0(0)
	mem[3] = 32'b10001100000010010000000000000100; //lw t1 4(0)
	mem[4] = 32'b10001100000010110000000000000000; //lw t3 0(0)
	
	
	//mem[2] = 32'b00000001000010011000000000100000; 
	//mem[3] = 32'b00000001000010011000100000100010; 
	//mem[4] = 32'b00000001000010011001000000100100; 
	//mem[5] = 32'b00000001000010011001100000100101; 
	//mem[6] = 32'b00000001000010011010000000101010;
	//mem[7] = 32'b00010010100000000000000000000110; 
	//mem[8] = 32'b00000001000010010101000000100000; 
	//mem[9] = 32'b00000001010010010101000000100000; 
	//mem[10] = 32'b00000001010010000101100000100000; 
	//mem[11] = 32'b10001100000101010000000000000100; 
	//mem[12] = 32'b00000001010101011011000000100000; 
	//mem[13] = 32'b00000010101010111011100000100000; 
	//mem[14] = 32'b10101100000101010000000000001000;
	//mem[15] = 32'b00001000000000000000000000000110;
	

	
end

always @(rdadd or reset) begin
	if (reset==1) begin
	
	mem[0] = 32'b00100000000010000000000000100000; //addi  t0 0 32
	mem[1] = 32'b00100000000010010000000000110111; //addi  t1 0 55
	mem[2] = 32'b10101100000010010000000000000000; //sw t1  0(0)
	mem[3] = 32'b10001100000010010000000000000100; //lw t1 4(0)
	mem[4] = 32'b10001100000010110000000000000000; //lw t3 0(0)
	
	
	end
	else begin
	add=rdadd/4;
	out=mem[add];
	end
end
endmodule
